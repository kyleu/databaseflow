general.ok = ok
general.loading = Läser in...
general.refresh = Uppdatera
general.cancel = Annullera
general.close = Stänga
general.previous = Tidigare
general.next = Nästa
general.coming.soon = Kommer snart
th.cancel = Annullera
th.column = Typ
th.columns = kolumner
th.connection = Förbindelse
th.cost = Kosta
th.default = Standard
th.definition = Definition
th.delete = Radera
th.description = Beskrivning
th.edit = Redigera
th.filter = Filtrera
th.foreign.keys = Utländska nycklar
th.indexes = index
th.name = namn
th.not.null = Inte Null
th.occurred = Inträffade
th.output = Produktion
th.owner = Ägare
th.parameters = parametrar
th.primary.key = Primärnyckel
th.properties = Egenskaper
th.read = Läsa
th.returns.result = Returnerar resultat
th.rows = rader
th.save = Spara
th.save.new = Spara som ny
th.settings = inställningar
th.source.columns = Källkolumner
th.sql = SQL
th.status = Status
th.target.columns = Målkolumner
th.target.table = Måltabell
th.title = Titel
th.type = Typ
th.unique = Unik
th.unknown = Okänd
history.title = Query History
history.remove.all = Ta bort hela historiken
history.no.records = Det verkar som om du inte har kört några frågor för den här databasen.
query.explain = Förklara
query.analyze = Analysera
query.export = Exportera
query.share = Dela med sig
query.chart = Diagram
query.data = Data
query.run = Springa
query.run.all = Kör alla
query.run.active = Kör Aktiv
query.run.selection = Kör markering
query.call = Samtalsproceduren
query.active.filter = Aktivt filter
query.no.rows.returned = Inga rader returnerade
query.insert = Lägg till ny rad
query.update = Uppdatera rad
query.insert.title = Ny [{0}] rad
query.update.title = Redigera [{0}] Rad ({1})
query.open.query = Ny fråga
query.view.first = Visa först 100 rader
query.load.more = Ladda {0} Fler rader
query.no.more.rows = Inga fler rader tillgängliga
query.plan = Query Plan
query.raw.plan = Visa Raw Plan
query.plan.estimated.rows = Est rader
query.error = Frågefel
query.plan.error = Planera fel
query.unsaved.changes = Den här frågan har inte sparat ändringar.
query.default.name = Ej sparad fråga {0}
query.open.relation = Öppna [{0}] med filter [{1}].
query.index.error = Ett fel uppstod vid index {0}.
query.chart.loading = Laddar diagramalternativ ...
feedback.title = Återkoppling
feedback.notice = Tack för din feedback.
feedback.email = E-postadress
feedback.prompt = Ange din feedback
feedback.submit = Skicka feedback
list.saved.queries = Sparade frågor
list.shared.results = Delade resultat
list.tables = tabeller
list.views = Visningar
list.procedures = Rutiner
list.this.connection = Den här anslutningen
list.unknown.connection = Okänd anslutning
list.all.connections = Alla anslutningar
list.filter = Filtrera {0}
graphql.title = GraphQL
help.title = {0} Hjälp
help.global.shortcuts = Globala genvägar
help.editor.shortcuts = Redigeringsgenvägar
help.tips.and.tricks = Tips och tricks
help.connection.status = Ansluten till servern med latens på [{0} ms].
help.hotkey.save.query = Spara fråga
help.hotkey.run.active.query = Kör aktiv fråga
help.hotkey.run.all.queries = Kör alla frågor
help.hotkey.leave.editor = Lämna redaktör
help.hotkey.help = Hjälpa
help.hotkey.search = Sök
help.hotkey.refresh.schema = Uppdatera schema
help.hotkey.new.query = Ny fråga
help.hotkey.focus.editor = Fokusera SQL Editor
help.hotkey.close.tab = Stäng fliken
help.hotkey.next.tab = Välj Nästa flik
help.hotkey.previous.tab = Välj Föregående flik
help.tip.theme = Du kan ändra färgschemat {0} från din profil när du är inloggad.
help.tip.hotkey.search = Tryck på [/] eller klicka i sökrutan för att börja filtrera databasobjekt.
help.tip.hotkey.new = Tryck på [+] när du är ute av en SQL-redigerare för att starta en ny fråga.
help.tip.hotkey.switch = Tryck på [eller] när utanför en SQL-redigerare för att växla mellan flikar.
help.tip.new.tab = Nästan alla länkar i {0} kan öppnas i nya webbläsarflikar för enkla jämförelser mellan sidor.