general.back.title = Tillbaka till anslutningslista
general.sql = SQL
general.error = Fel
general.about = Handla om
general.save = Spara
general.cancel = Annullera
general.loading = Läser in...
general.delete = Radera
general.ok = ok
general.edit = Redigera
th.columns = Cols
th.connection = Förbindelse
th.created = Skapad
th.duration = Dur
th.edition = Utgåva
th.elapsed = förfluten
th.email = E-post
th.export = Exportera
th.first = 1:a
th.import = Importera
th.issued = Utfärdad
th.last.accessed = Senast åtkomlig
th.name = namn
th.occurred = Inträffade
th.owner = Ägare
th.role = Roll
th.rows = rader
th.status = Status
th.table = Tabell
th.theme = Tema
th.type = Typ
th.username = Användarnamn
index.no.connections = Lägg till din första anslutning genom att klicka på länken nedan.
index.new.connection = Ny anslutning
registration.title = Registrera
registration.call.to.action = Registrera dig för {0}
registration.notice = Du skapar ett konto för den här lokala installationen av {0}. 
registration.register = Bli Medlem
registration.email.taken = Den e-postadressen används redan
registration.form.username = namn
registration.form.email = E-postadress
registration.form.password = Lösenord
registration.form.password.confirm = Bekräfta lösenord
registration.passwords.do.not.match = Lösenorden matchar inte
registration.already.member = redan medlem?
registration.disabled = Du kan inte registrera dig just nu. 
authentication.call.to.action = Logga in på {0}
authentication.notice = Detta konto är endast för denna installation av {0}. 
authentication.sign.in = Logga in
authentication.sign.out = Logga ut
authentication.form.email = E-postadress
authentication.form.password = Lösenord
authentication.invalid.credentials = Ogiltiga uppgifter
authentication.not.member = Inte en medlem?
authentication.registration.disabled = Registrering är inaktiverad på den här servern. 
profile.title = Profil
profile.save = Spara ändringar
profile.cancel = Annullera
profile.change.password = Ändra lösenord
profile.change.password.old = Gammalt lösenord
profile.change.password.new = nytt lösenord
profile.change.password.confirm = Bekräfta nytt lösenord
profile.form.username = Användarnamn
profile.form.language = Språk
profile.form.theme = Tema
activity.title = Aktivitet
activity.profile.title = Användaraktivitet
activity.admin.title = Systemaktivitet
activity.no.results = Ingen aktivitet registrerad i databasen.
activity.load.more = Ladda {0} Mer
activity.remove.confirm = Borttagen aktivitet [{0}]
activity.remove.all = Ta bort all aktivitet
activity.remove.ok = Ta bort aktivitet [{0}].
activity.remove.all.confirm = Ta bort all systemaktivitet.
activity.remove.all.user.confirm = Ta bort all användaraktivitet.
activity.confirm.remove.user = Är du säker på att du vill ta bort all din verksamhet?
activity.confirm.remove.all = Är du säker på att du vill ha all aktivitet från systemet?
permissions.everyone = Alla
permissions.registered.users = registrerade användare
permissions.administrators = Administratörer
permissions.only.myself = Bara mig själv
permissions.visitor.text = Av alla
permissions.user.text = Av alla registrerade användare
permissions.administrators.text = Av administratörer
permissions.private.text = Bara av dig
connection.permissions.available.to = Tillgänglig för
connection.permissions.editable.by = Redigerbar av
connection.name = Anslutningsnamn
connection.engine = Databasmotor
connection.username = Användarnamn
connection.password = Lösenord
connection.url = URL
connection.fields = Fields
connection.host = Värd
connection.port = Hamn
connection.db.name = Databas namn
connection.jdbc.url = Jdbc URL
connection.description = Beskrivning
connection.new.title = Ny anslutning
connection.permission.denied = Du har inte behörighet att lägga till en databasanslutning.
query.title = Fråga
query.loading = Laddar {0} ...
query.search = Sök
query.tx.begin = Börja Transaktion
query.tx.none = Ingen aktiv transaktion.
query.tx.commit = Commit Transaction
query.tx.rollback = Rulla tillbaka
query.sidenav.loading = Läser in...
query.sidenav.new = Ny fråga
query.sidenav.history = Query History
query.sidenav.refresh = Uppdatera schema
query.sidenav.saved.queries = Sparade frågor
query.sidenav.shared.results = Delade resultat
query.sidenav.tables = tabeller
query.sidenav.views = Visningar
query.sidenav.procedures = Lagrade procedurer
query.sidenav.graphql = GraphQL
query.sidenav.help = Hjälpa
query.sidenav.feedback = Återkoppling
query.sidenav.about = Om {0}
query.share = Dela med sig
query.insert = Sätt in rad
query.edit = Redigera
result.remove.confirm = Raderat resultat [{0}].
result.remove.orphan = Ta bort föräldralösa bord [{0}].
shared.results.title = Delade resultat
shared.results.personal.title = Mina delade resultat
shared.results.public.title = Public Shared Results
shared.results.public.none = Inga offentliga delade resultat tillgängliga.
graphql.title = GraphQL
socket.connect.error = Ett fel försökte ansluta till databasen.
socket.connect.failed = Anslutningen misslyckades
socket.too.many.users = Personal Edition tillåter endast en användare att ansluta åt gången och [{0}] är redan ansluten.
socket.duplicate.transaction = Redan i en transaktion.
socket.no.transaction = För närvarande inte i en transaktion.
modal.confirm.prompt = Är du säker?
modal.export.action = Exportera
modal.export.csv = Kommaseparerade värden
modal.export.excel = Microsoft excel
modal.reconnect.prompt = Anslutningsfel. 
modal.reconnect.action = Anslut
modal.save.query.name = Fråga namn
modal.save.description = Beskrivning
modal.save.available.from = Tillgänglig från
modal.save.all.databases = Alla databaser
modal.save.this.database = Endast denna databas
modal.share.results.title = Titel
modal.share.results.description = Beskrivning
user.password.changed = Lösenordet ändrat.
user.password.check.fail = Gammalt lösenord matchar inte ({0}).
admin.title = inställningar
admin.back.title = Tillbaka
admin.index.title = {0} Administration
admin.index.prompt = Använd menyn ovan eller länkarna nedan för att komma igång!
admin.status.link = Status
admin.status.title = {0} Status
admin.status.description = Visa systemstatus.
admin.status.metrics.title = System Metrics
admin.status.file.loaded = Laddad från {0}
admin.status.db.loaded = {0} databas, laddad från {1}
admin.settings.link = Inställningar
admin.settings.title = Systeminställningar
admin.settings.description = Redigera systeminställningar.
admin.settings.invalid = Försök att spara ogiltig inställning [{0}].
admin.users.link = användare
admin.users.title = Användarhantering
admin.users.description = Hantera systemets användare.
admin.results.link = Resultat
admin.results.title = Cached Query Results
admin.results.description = Visa cachelagrade sökresultat som har sparats.
admin.activity.link = Aktivitet
admin.activity.title = Användaraktivitet
admin.activity.description = Visa systemaktiviteten för alla användare i systemet.
admin.users.new = Ny användare
admin.users.confirm = Är du säker på att du vill radera den här användaren ({0})?
error.admin.required = Du måste ha administratörsrättigheter för att komma åt den sidan.
error.not.logged.in = På något sätt inte inloggad.
error.must.sign.in = Du måste logga in eller registrera innan du öppnar {0}.
error.missing.parameter = Saknar [{0}] parameter.
error.unknown.format = Okänt format [{0}].
error.exception.encountered = Det gick inte att exportera fråga: [{0}: {1}].
error.sign.in.disabled = Endast administratörer kan logga in just nu. 
error.missing.user = Det gick inte att hitta användaren {0}.
error.cannot.sign.up = Det gick inte att registrera sig vid denna tidpunkt. 
error.empty = {0} krävs.
error.invalid.user = Ogiltig användare [{0}].
error.remove.self = Du kan inte ta bort din egen administratörsroll.