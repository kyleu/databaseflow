general.save = Spara
general.about = Om
th.email = E-post
th.name = Namn
index.splash = Vi arbetar hårt på en ny idé. Kommer snart!
index.features.link = Funktioner
index.download.link = Ladda ner
index.versions.link = Versioner
index.admin.link = Admin
index.welcome1 = {0} är det bästa sättet att fråga och rapport på din egen data.
index.welcome2 = Du kan köra {0} lokalt för eget bruk, eller installera till en gemensam server för hela laget.
downloads.title = Nedladdningar
platform.osx = macOS
platform.windows = Windows
platform.linux = Linux
platform.docker = Docker
license.title = Få en Licens
license.personal = Få En Gratis Personlig Edition-Licens
license.team = Köp Team Edition Nu
features.a = Sparade frågor
features.b = Redaktör för komplettera automatiskt
features.c = Gränssnitt
features.d = Detaljer av tabeller, vyer och procedurer
features.e = Länka till relaterade tabeller
features.f = Behörigheter för databaser och frågor
features.g = Material och design
features.h = Responsiv design med mobilt stöd
features.i = Stöder H2, MySQL, Oracle, PostgreSQL, och SQL Server
features.j = Lokalt installerade program
features.k = Inga annonser, spår eller webbplatser från tredje part
features.l = Visa kolumner, index, nyckel
newsletter.title = Nyhetsbrev
newsletter.subscribe = Prenumerera
feedback.title = Feedback
feedback.action = Lämna Feedback
feedback.email = E-Postadress
feedback.submit = Skicka Feedback
license.download = Ladda Ner Licensfil
license.copy = Kopiera Licens till Urklipp
license.success = Din {0} Licens
license.continue = Fortsätt
license.form.name = Namn
license.form.email = E-post
license.form.prompt = Fyll i denna blankett, och du kommer att få din licens omedelbart.
license.form.personal = Ny Personlig Licens
purchase.title = Köp Licens
static.copyright = © 2016 {0}