general.save = Spara
general.about = Om
general.back = Tillbaka
th.email = E-post
th.name = Namn
index.splash = Vi arbetar hårt på en ny idé. Kommer snart!
index.features.link = Funktioner
index.demo.link = Visa Demo
index.download.link = Ladda ner
index.admin.link = Admin
index.welcome1 = Det bästa sättet att fråga och rapport på din egen data.
index.welcome2 = Du kan köra {0} lokalt för eget bruk, eller installera till en gemensam server för hela laget.
index.hero.title = Det bästa sättet att fråga och visualisera din databas.
index.hero.subtitle1 = {0} är en egen värd samarbete SQL-klient och kartläggning program som fungerar med din databas.
index.hero.subtitle2 = Du kan köra {0} lokalt för eget bruk, eller installera till en gemensam server för hela laget.
downloads.title = Nedladdningar
downloads.hero.title = Komma igång med {0} direkt.
downloads.hero.subtitle1 = Nedladdningar som är tillgängliga för alla större plattformar.
platform.osx = macOS
platform.windows = Windows
platform.linux = Linux
platform.docker = Docker
platform.universal = Universal (kräver Java 8)
newsletter.title = Nyhetsbrev
newsletter.subscribe = Prenumerera
feedback.title = Feedback
feedback.action = Lämna Feedback
feedback.email = E-Postadress
feedback.submit = Skicka Feedback
versions.hero.title = Välj den version som är rätt för dig.
versions.hero.subtitle1 = Prova {0} under trettio dagar, eller köpa en licens för dig själv eller hela laget.
features.hero.title = {0} är en modern webb-baserade SQL-klient.
features.hero.subtitle1 = Med hjälp av streaming webb-teknik, {0} hjälper dig att komma åt dina data från valfri enhet.
technology.hero.title = {0} bygger på enorma projekt med öppen källkod.
technology.hero.subtitle1 = Här är några av dem.
database.hero.title = {0} är den bästa SQL-klient för att arbeta med {1}
database.postgresql.subtitle = {1} är vår primära stöd databas, vi stöd för normala installationer, Amazon RDS eller Rödförskjutning, och Greenplum.
purchase.title = Köp {0} Edition-Licens
footer.newsletter = Nyhetsbrev
footer.technology = Teknik
footer.feedback = Feedback
