general.save = Spara
general.about = Handla om
general.back = Tillbaka
th.email = E-post
th.name = namn
index.splash = Vi arbetar hårt med en ny idé. 
index.features.link = Funktioner
index.demo.link = Visa demo
index.download.link = Ladda ner
index.admin.link = Administration
index.welcome1 = Det bästa sättet att fråga och rapportera om dina egna data.
index.welcome2 = Du kan köra {0} lokalt för egen användning, eller installera till en gemensam server för hela laget.
index.hero.title = Det bästa sättet att fråga och visualisera din databas.
index.hero.subtitle1 = {0} är en självhävd samverkande SQL-klient och kartläggningsprogram som fungerar med din databas.
index.hero.subtitle2 = Du kan köra {0} lokalt för egen användning, eller installera till en gemensam server för hela laget.
github.title = github
downloads.title = Ladda ner nu
downloads.hero.title = Kom igång med {0} direkt.
downloads.hero.subtitle1 = Fri programvara, ingen registrering krävs. 
platform.osx = Mac OS
platform.windows = Windows
platform.linux = Linux
platform.docker = Hamnarbetare
platform.universal = Universal (kräver Java 8)
newsletter.title = Nyhetsbrev
newsletter.subscribe = Prenumerera
feedback.title = Återkoppling
feedback.action = Lämna feedback
feedback.email = E-postadress
feedback.submit = Skicka feedback
features.hero.title = {0} är en modern webbaserad SQL-klient.
features.hero.subtitle1 = Med hjälp av strömmande webbteknik hjälper {0} dig åt dig åtkomst till dina data från vilken enhet som helst.
technology.hero.title = {0} bygger på enorma open source-projekt.
technology.hero.subtitle1 = Här är några av dem.
database.hero.title = {0} är den bästa SQL-klienten för att arbeta med {1}
database.postgresql.subtitle = {0} är vår primära databas, vi stöder normala installationer, Amazon RDS eller Redshift och Greenplum.
footer.newsletter = Nyhetsbrev
footer.technology = Teknologi
footer.feedback = Återkoppling