general.back.title = Tillbaka till Anslutning Lista
general.sql = SQL
general.error = Fel
general.about = Om
general.save = Spara
general.cancel = Avbryt
general.delete = Ta bort
general.ok = OK
general.edit = Ändra
th.columns = Cols
th.connection = Anslutning
th.created = Skapad
th.duration = Dur
th.edition = Edition
th.elapsed = Uppspelad
th.email = E-post
th.export = Export
th.first = 1: a
th.import = Importera
th.issued = Utfärdat
th.last.accessed = Senast Öppnad
th.name = Namn
th.occurred = Inträffade
th.owner = Ägare
th.role = Roll
th.rows = Rader
th.status = Status
th.table = Tabell
th.theme = Tema
th.type = Typ
th.username = Användarnamn
index.welcome = Välkommen till {0}! Här"sa några ord om appen. Kanske en slogan eller något.
index.no.connections = Lägg till din första anslutningen genom att klicka på länken nedan.
index.new.connection = Ny Anslutning
license.new.form = Licens Detaljer
license.paste = Klistra in din licens i formuläret nedan.
license.missing = Saknas licens innehåll.
license.success = Licens uppdaterats.
registration.title = Registrera dig
registration.call.to.action = Registrera dig för {0}
registration.register = Registrera Dig
registration.email.taken = E-postadressen används redan
registration.form.username = Namn
registration.form.email = E-Postadress
registration.form.password = Lösenord
registration.form.password.confirm = Bekräfta Lösenord
registration.passwords.do.not.match = Lösenorden matchar inte
registration.already.member = Är du redan medlem?
registration.disabled = Du kan inte anmäla dig vid denna tid. Kontakta din administratör.
authentication.call.to.action = Logga in på {0}
authentication.sign.in = Logga In
authentication.sign.out = Logga Ut
authentication.form.email = E-Postadress
authentication.form.password = Lösenord
authentication.invalid.credentials = Ogiltiga referenser
authentication.not.member = Inte medlem?
authentication.registration.disabled = Registrering är inaktiverad på servern. Kontakta din administratör för att få ett konto.
profile.title = Profil
profile.save = Spara Ändringar
profile.cancel = Avbryt
profile.change.password = Ändra Lösenord
profile.change.password.old = Gammalt Lösenord
profile.change.password.new = Nytt Lösenord
profile.change.password.confirm = Bekräfta Nytt Lösenord
profile.form.username = Användarnamn
profile.form.language = Språk
profile.form.theme = Tema
activity.title = Aktivitet
activity.profile.title = Användarens Aktivitet
activity.admin.title = Systemet Aktivitet
activity.no.results = Ingen aktivitet registreras i databasen.
activity.load.more = Ladda {0} Mer
activity.remove.confirm = Bort aktivitet [{0}]
activity.remove.all = Ta Bort All Aktivitet
activity.remove.ok = Bort aktivitet [{0}].
activity.remove.all.confirm = Tagit bort alla system för aktivitet.
activity.remove.all.user.confirm = Bort all användaraktivitet.
activity.confirm.remove.user = Är du säker på att du vill ta bort alla dina aktiviteter?
activity.confirm.remove.all = Är du säker på att du vill att all aktivitet från systemet?
permissions.everyone = Alla
permissions.registered.users = Registrerade Användare
permissions.administrators = Administratörer
permissions.only.myself = Bara Mig Själv
permissions.visitor.text = alla
permissions.user.text = alla registrerade användare
permissions.administrators.text = administratörer
permissions.only.myself.text = bara du
connection.permissions.available.to = Tillgänglig För
connection.permissions.editable.by = Redigeras Av
connection.name = Anslutningsnamn
connection.engine = Databasmotorn
connection.username = Användarnamn
connection.password = Lösenord
connection.url = URL
connection.fields = Fält
connection.host = Värd
connection.port = Port
connection.db.name = Databas Namn
connection.jdbc.url = Jdbc-URL
connection.description = Beskrivning
connection.new.title = Ny Anslutning
connection.permission.denied = Du har inte behörighet att lägga till en koppling till en databas.
query.title = Fråga
query.loading = Fylla på {0}...
query.search = Sök
query.tx.begin = Börja Transaktion
query.tx.none = Ingen aktiv transaktion.
query.tx.commit = Begå Transaktion
query.tx.rollback = Rollback
query.sidenav.loading = Laddar...
query.sidenav.new = Ny Fråga
query.sidenav.history = Frågan Historia
query.sidenav.refresh = Uppdatera Schema
query.sidenav.saved.queries = Sparade Frågor
query.sidenav.shared.results = Gemensamt Resultat
query.sidenav.tables = Tabeller
query.sidenav.views = Visningar
query.sidenav.procedures = Lagrade Procedurer
query.sidenav.help = Hjälp
query.sidenav.feedback = Feedback
query.sidenav.about = Om {0}
query.share = Dela
result.remove.confirm = Bort resultat [{0}].
result.remove.orphan = Ta bort anonyma bord [{0}].
shared.results.title = Gemensamt Resultat
shared.results.personal.title = Mina Delade Resultat
shared.results.public.title = Allmänna Gemensamt Resultat
shared.results.public.none = Inga offentliga gemensamt resultat.
socket.connect.error = Fel vid försök att ansluta till databasen.
socket.connect.failed = Anslutning Misslyckades
socket.too.many.users = Personal Edition endast tillåter en användare att ansluta på en gång, och [{0}] är redan ansluten.
socket.duplicate.transaction = Redan i en transaktion.
socket.no.transaction = För närvarande inte i en transaktion.
modal.confirm.prompt = Är du säker?
modal.export.action = Export
modal.export.csv = Kommaavgränsade Värden
modal.export.excel = Microsoft Excel
modal.reconnect.prompt = Anslutningsfel. Vill du försöka igen?
modal.reconnect.action = Återanslut
modal.save.query.name = Fråga Namn
modal.save.description = Beskrivning
modal.save.available.from = Tillgängligt Från
modal.save.all.databases = Alla Databaser
modal.save.this.database = Denna Databas Endast
modal.share.results.title = Titel
modal.share.results.description = Beskrivning
user.password.changed = Lösenord ändrat.
user.password.check.fail = Gamla lösenordet matchar inte ({0}).
admin.title = Administration
admin.index.title = {0} Administration
admin.index.prompt = Använd menyn ovan eller länkarna nedan för att komma igång!
admin.settings.link = Inställningar
admin.settings.title = System Inställningar
admin.settings.description = Redigera system inställningar och preferenser.
admin.settings.invalid = Försök att spara ogiltiga inställningen [{0}].
admin.users.link = Användare
admin.users.title = Användarhantering
admin.users.description = Hantera användare av systemet.
admin.results.link = Resultat
admin.results.title = Cachade Frågeresultat
admin.results.description = Visa cachade fråga resultaten att ha sparats.
admin.activity.link = Aktivitet
admin.activity.title = Användarens Aktivitet
admin.activity.description = Visa system aktivitet för alla användare i systemet.
admin.users.new = Ny Användare
admin.users.confirm = Är du säker på att du vill ta bort den här användaren ({0})?
error.admin.required = Du måste ha administratörsbehörighet för att komma åt sidan.
error.not.logged.in = På något sätt inte är inloggad.
error.must.sign.in = Du måste logga in eller registrera dig innan du får åtkomst till {0}.
error.missing.parameter = Saknas [{0}] parameter.
error.unknown.format = Okänt format [{0}].
error.exception.encountered = Det går inte att exportera fråga: [{0}: {1}].
error.missing.user = Kunde inte hitta användaren {0}.
error.cannot.sign.up = Det går inte att logga upp vid den här tiden. Kontakta din administratör.
error.empty = {0} är som krävs.
error.invalid.user = Ogiltig användare [{0}].
error.remove.self = Du kan inte ta bort dina egna rollen admin.
static.copyright = © 2016 {0}