general.save = Spara
general.about = Handla om
general.back = Tillbaka
th.email = E-post
th.name = namn
index.splash = Vi arbetar hårt med en ny idé.
index.features.link = Funktioner
index.demo.link = Visa demo
index.download.link = Ladda ner
index.github.link = github
index.admin.link = Administration
index.hero.title = Fråga din databas med ett modernt webbgränssnitt för SQL och GraphQL.
index.hero.subtitle1 = {0} är en öppen källkod, självhävd SQL-klient, GraphQL-server och kartläggningsprogram som fungerar med din databas.
index.hero.subtitle2 = Visualisera scheman, frågeplaner, diagram och resultat.
downloads.title = Ladda ner nu
downloads.hero.title = Kom igång med {0} direkt.
downloads.hero.subtitle1 = Gratis programvara, ingen registrering krävs.
downloads.dependency.java8 = Java 8 krävs
features.manage.title = Hantera dina data
features.manage.content = Kör SQL-frågor, utforska databasobjekt och dela och visualisera resultaten.
features.editor.title = Avancerad SQL Editor
features.editor.content = Syntaxutmärkning och automatisk slutförande gör det enkelt att skriva komplicerade frågor.
features.charting.title = kartläggning
features.charting.content = Vi använder plotly.js för att få dig de bästa kartorna tillgängliga.
features.plan.title = Query Plan
features.plan.content = Visualisera resultatet av dina frågor med en sofistikerad planvisare.
features.graphql.title = GraphQL
features.graphql.content = Använd GraphQLs kraft för att utforska och upptäcka din databas.
features.schema.title = Utforska ditt schema
features.schema.content = Visualisera relationer och kolumner i ditt databasschema.
features.responsive.title = Responsive Interface
features.responsive.content = High Definition näthinnans grafik och ett lyhörd gränssnitt hjälper dig att navigera dina data på vilken enhet som helst.
features.databases.title = Databasstöd
features.databases.content = Database Flow stöder de mest populära databasmotorerna och ger funktioner som hjälper dig att få ut mesta möjliga av dina data.
features.filter.title = Resultatfiltrering
features.filter.content = Sortera och filtrera dina resultat utan att köra din fråga igen.
features.history.title = Query History
features.history.content = Frågehistorik och revisionsloggar ser till att du aldrig glömmer de frågor du skriver.
newsletter.title = Nyhetsbrev
newsletter.subscribe = Prenumerera
feedback.title = Återkoppling
feedback.action = Lämna feedback
feedback.email = E-postadress
feedback.submit = Skicka feedback
features.hero.title = {0} är en modern webbaserad SQL-klient och GraphQL-server.
features.hero.subtitle1 = Med hjälp av strömmande webbteknik hjälper {0} dig åt dig åtkomst till dina data från vilken enhet som helst.
technology.hero.title = {0} bygger på enorma open source-projekt.
technology.hero.subtitle1 = Här är några av dem.
database.supported.databases = Stödda databaser
database.hero.title = {0} är en egen värd SQL-klient och GraphQL sever för att arbeta med {1}.
database.db2.subtitle = Vi har testat grundläggande funktionalitet för {0}.
database.h2.subtitle = Fråga och visualisera dina {0} databaser med SQL eller GraphQL.
database.informix.subtitle = Vi har testat grundläggande funktionalitet för {0}.
database.mysql.subtitle = Fråga och visualisera dina {0} databaser och fråga planer, med hjälp av SQL eller GraphQL.
database.oracle.subtitle = Vi har testat grundläggande funktionalitet för {0}.
database.postgresql.subtitle = {0} är vår primära databas, vi stöder normala installationer, Amazon RDS eller Redshift och Greenplum.
database.sqlite.subtitle = Fråga och visualisera dina {0} databaser och fråga planer, med hjälp av SQL eller GraphQL.
database.sqlserver.subtitle = Vi har testat grundläggande funktionalitet för {0}.
footer.newsletter = Nyhetsbrev
footer.technology = Teknologi
footer.feedback = Återkoppling