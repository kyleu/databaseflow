general.ok = OK
general.loading = Laddar...
general.refresh = Uppdatera
general.cancel = Avbryt
general.close = Stäng
general.previous = Föregående
general.next = Nästa
general.coming.soon = Kommer Snart
th.cancel = Avbryt
th.column = Typ
th.columns = Kolumner
th.connection = Anslutning
th.cost = Kostnad
th.default = Standard
th.definition = Definition
th.delete = Ta bort
th.description = Beskrivning
th.edit = Ändra
th.filter = Filter
th.foreign.keys = Främmande Nycklar
th.indexes = Index
th.name = Namn
th.not.null = Null
th.occurred = Inträffade
th.output = Utgång
th.owner = Ägare
th.parameters = Parametrar
th.primary.key = Primär Nyckel
th.properties = Egenskaper
th.read = Läs
th.returns.result = Returnerar Resultatet
th.rows = Rader
th.save = Spara
th.save.new = Spara som Ny
th.settings = Inställningar
th.source.columns = Källa Kolumner
th.sql = SQL
th.status = Status
th.target.columns = Målet Kolumner
th.target.table = Målet Tabellen
th.title = Titel
th.type = Typ
th.unique = Unik
th.unknown = Okänd
history.title = Frågan Historia
history.remove.all = Ta Bort All Historik
history.no.records = Det ser ut som att du inte köra alla frågor för den här databasen. Komma igång!
query.explain = Förklara
query.analyze = Analysera
query.export = Export
query.share = Dela
query.chart = Diagram
query.data = Data
query.run = Kör
query.run.all = Kör Alla
query.run.active = Kör Aktiv
query.run.selection = Kör Urval
query.call = Samtal Förfarande
query.active.filter = Aktiva Filter
query.no.rows.returned = Några rader tillbaka
query.insert = Lägg Till Ny Rad
query.view.first = Visa Första 100 Rader
query.load.more = Ladda {0} Fler Rader
query.no.more.rows = Inga fler rader finns
query.plan = Fråga Plan
query.raw.plan = Visa Raw-Plan
query.plan.estimated.rows = Est Rader
query.error = Frågan Fel
query.plan.error = Plan För Fel
query.unsaved.changes = Denna fråga har osparade ändringar.
query.default.name = Osparade Frågan {0}
query.open.relation = Öppna [{0}] tabell filtreras där [{1}].
query.index.error = Fel som uppstått på index {0}.
query.chart.loading = Laddar diagram alternativ...
feedback.title = Feedback
feedback.notice = Tack för din feedback. Detta kommer att skicka ditt meddelande direkt till skaparna av {0}. Om du vill bli meddelad när vi svarar, vänligen inkludera en e-postadress.
feedback.email = E-Postadress
feedback.prompt = Skriv in din feedback
feedback.submit = Lämna Feedback
list.saved.queries = Sparade Frågor
list.shared.results = Gemensamt Resultat
list.tables = Tabeller
list.views = Visningar
list.procedures = Förfaranden
list.this.connection = Denna Anslutning
list.unknown.connection = Okänd Anslutning
list.all.connections = Alla Anslutningar
list.filter = Filtrera {0}
help.title = {0} Hjälp
help.global.shortcuts = Globala Genvägar
help.editor.shortcuts = Redaktör Genvägar
help.tips.and.tricks = Tips och Tricks
help.connection.status = Ansluten med en latens på [{0}ms]. Vi har skickat {1} och fick {2} meddelanden.
help.hotkey.save.query = Spara Sökning
help.hotkey.run.active.query = Kör Aktivt Fråga
help.hotkey.run.all.queries = Kör Alla Frågor
help.hotkey.leave.editor = Lämna Redaktör
help.hotkey.help = Hjälp
help.hotkey.search = Sök
help.hotkey.refresh.schema = Uppdatera Schema
help.hotkey.new.query = Ny Fråga
help.hotkey.focus.editor = Fokus SQL-Editor
help.hotkey.close.tab = Stäng Flik
help.hotkey.next.tab = Välj Nästa Flik
help.hotkey.previous.tab = Välj Föregående Flik
help.tip.theme = Du kan ändra färgschemat för {0} från din profil när du är inloggad.
help.tip.hotkey.search = Tryck på [/] eller klicka i rutan sök för att starta filtrering av databas-objekt.
help.tip.hotkey.new = Tryck på [+] när du befinner dig utanför i en sql-editor för att starta en ny sökning.
help.tip.hotkey.switch = Tryck på [] när du är utanför av en sql-editor för att växla mellan flikarna.
help.tip.new.tab = Nästan alla länkar i {0} kan öppnas i nya flikar i webbläsaren för enkel sida vid sida jämförelser.