general.save = Spara
general.about = Om
th.email = E-post
th.name = Namn
index.splash = Vi arbetar hårt på en ny idé. Kommer snart!
index.features.link = Funktioner
index.download.link = Ladda ner
index.versions.link = Versioner
index.admin.link = Admin
downloads.title = Nedladdningar
platform.osx = macOS
platform.windows = Windows
platform.linux = Linux
platform.docker = Docker
license.title = Få en Licens
license.personal = Få En Gratis Personlig Edition-Licens
license.team = Köp Team Edition Nu
newsletter.title = Nyhetsbrev
newsletter.subscribe = Prenumerera
feedback.title = Feedback
feedback.action = Lämna Feedback
feedback.email = E-Postadress
feedback.submit = Skicka Feedback
license.download = Ladda Ner Licensfil
license.copy = Kopiera Licens till Urklipp
license.success = Din Databas Flöde Licens
license.continue = Fortsätt
license.form.name = Namn
license.form.email = E-post
license.form.prompt = Fyll i denna blankett, och du kommer att få din licens omedelbart.
license.form.personal = Ny Personlig Licens
purchase.description = Fyll i denna blankett, och du kommer att få din licens omedelbart.
purchase.title = Köp Licens
static.copyright = © 2016 {0}